-- megafunction wizard: %ALTMULT_ADD%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: ALTMULT_ADD 

-- ============================================================
-- File Name: altmult_add0.vhd
-- Megafunction Name(s):
-- 			ALTMULT_ADD
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 304 01/25/2010 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2010 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY altmult_add0 IS
	PORT
	(
		dataa_0		: IN STD_LOGIC_VECTOR (15 DOWNTO 0) :=  (OTHERS => '0');
		datab_0		: IN STD_LOGIC_VECTOR (15 DOWNTO 0) :=  (OTHERS => '0');
		result		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
END altmult_add0;


ARCHITECTURE SYN OF altmult_add0 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (15 DOWNTO 0);



	COMPONENT altmult_add
	GENERIC (
		addnsub_multiplier_pipeline_register1		: STRING;
		addnsub_multiplier_register1		: STRING;
		dedicated_multiplier_circuitry		: STRING;
		input_register_a0		: STRING;
		input_register_b0		: STRING;
		input_source_a0		: STRING;
		input_source_b0		: STRING;
		intended_device_family		: STRING;
		lpm_type		: STRING;
		multiplier1_direction		: STRING;
		multiplier_register0		: STRING;
		number_of_multipliers		: NATURAL;
		output_register		: STRING;
		port_addnsub1		: STRING;
		port_signa		: STRING;
		port_signb		: STRING;
		representation_a		: STRING;
		representation_b		: STRING;
		signed_pipeline_register_a		: STRING;
		signed_pipeline_register_b		: STRING;
		signed_register_a		: STRING;
		signed_register_b		: STRING;
		width_a		: NATURAL;
		width_b		: NATURAL;
		width_result		: NATURAL
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(15 DOWNTO 0);

	ALTMULT_ADD_component : ALTMULT_ADD
	GENERIC MAP (
		addnsub_multiplier_pipeline_register1 => "UNREGISTERED",
		addnsub_multiplier_register1 => "UNREGISTERED",
		dedicated_multiplier_circuitry => "AUTO",
		input_register_a0 => "UNREGISTERED",
		input_register_b0 => "UNREGISTERED",
		input_source_a0 => "DATAA",
		input_source_b0 => "DATAB",
		intended_device_family => "Cyclone III",
		lpm_type => "altmult_add",
		multiplier1_direction => "ADD",
		multiplier_register0 => "UNREGISTERED",
		number_of_multipliers => 1,
		output_register => "UNREGISTERED",
		port_addnsub1 => "PORT_UNUSED",
		port_signa => "PORT_UNUSED",
		port_signb => "PORT_UNUSED",
		representation_a => "SIGNED",
		representation_b => "SIGNED",
		signed_pipeline_register_a => "UNREGISTERED",
		signed_pipeline_register_b => "UNREGISTERED",
		signed_register_a => "UNREGISTERED",
		signed_register_b => "UNREGISTERED",
		width_a => 16,
		width_b => 16,
		width_result => 16
	)
	PORT MAP (
		dataa => dataa_0,
		datab => datab_0,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADDER1_ROUND_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER1_ROUND_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER1_ROUND_OP STRING "Enabled"
-- Retrieval info: PRIVATE: ADDER1_ROUND_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER1_ROUND_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER1_ROUND_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: ADDER1_ROUND_REG STRING "0"
-- Retrieval info: PRIVATE: ADDER1_SAT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER1_SAT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER1_SAT_OP STRING "Enabled"
-- Retrieval info: PRIVATE: ADDER1_SAT_OVERFLOW_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER1_SAT_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER1_SAT_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER1_SAT_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: ADDER1_SAT_REG STRING "0"
-- Retrieval info: PRIVATE: ADDER3_ROUND_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER3_ROUND_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER3_ROUND_OP STRING "Enabled"
-- Retrieval info: PRIVATE: ADDER3_ROUND_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDER3_ROUND_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDER3_ROUND_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: ADDER3_ROUND_REG STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB1_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB1_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB1_REG STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB3_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: ADDNSUB3_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: ADDNSUB3_REG STRING "0"
-- Retrieval info: PRIVATE: ADD_ENABLE NUMERIC "0"
-- Retrieval info: PRIVATE: ALL_REG_ACLR NUMERIC "0"
-- Retrieval info: PRIVATE: A_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: A_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: B_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: B_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: HAS_MAC STRING "0"
-- Retrieval info: PRIVATE: HAS_SAT_ROUND STRING "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEDICATED NUMERIC "0"
-- Retrieval info: PRIVATE: IMPL_STYLE_DEFAULT NUMERIC "1"
-- Retrieval info: PRIVATE: IMPL_STYLE_LCELL NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: MULT01_ROUND_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT01_ROUND_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT01_ROUND_OP STRING "Enabled"
-- Retrieval info: PRIVATE: MULT01_ROUND_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT01_ROUND_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT01_ROUND_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: MULT01_ROUND_REG STRING "0"
-- Retrieval info: PRIVATE: MULT01_SAT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT01_SAT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT01_SAT_OP STRING "Enabled"
-- Retrieval info: PRIVATE: MULT01_SAT_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT01_SAT_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT01_SAT_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: MULT01_SAT_REG STRING "0"
-- Retrieval info: PRIVATE: MULT0_SAT_OVERFLOW_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: MULT1_SAT_OVERFLOW_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: MULT23_ROUND_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT23_ROUND_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT23_ROUND_OP STRING "Enabled"
-- Retrieval info: PRIVATE: MULT23_ROUND_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT23_ROUND_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT23_ROUND_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: MULT23_ROUND_REG STRING "0"
-- Retrieval info: PRIVATE: MULT23_SAT_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT23_SAT_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT23_SAT_OP STRING "Enabled"
-- Retrieval info: PRIVATE: MULT23_SAT_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: MULT23_SAT_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: MULT23_SAT_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: MULT23_SAT_REG STRING "0"
-- Retrieval info: PRIVATE: MULT2_SAT_OVERFLOW_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: MULT3_SAT_OVERFLOW_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGA0 NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGB0 NUMERIC "0"
-- Retrieval info: PRIVATE: MULT_REGOUT0 NUMERIC "0"
-- Retrieval info: PRIVATE: NUM_MULT STRING "1"
-- Retrieval info: PRIVATE: OP1 STRING "Add"
-- Retrieval info: PRIVATE: OP3 STRING "Add"
-- Retrieval info: PRIVATE: OUTPUT_EXTRA_LAT NUMERIC "0"
-- Retrieval info: PRIVATE: OUTPUT_REG_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: OUTPUT_REG_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: Q_ACLR_SRC_MULT0 NUMERIC "3"
-- Retrieval info: PRIVATE: Q_CLK_SRC_MULT0 NUMERIC "0"
-- Retrieval info: PRIVATE: REG_OUT NUMERIC "0"
-- Retrieval info: PRIVATE: RNFORMAT STRING "16"
-- Retrieval info: PRIVATE: RQFORMAT STRING "Q1.15"
-- Retrieval info: PRIVATE: RTS_WIDTH STRING "16"
-- Retrieval info: PRIVATE: SAME_CONFIG NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_A0 NUMERIC "1"
-- Retrieval info: PRIVATE: SAME_CONTROL_SRC_B0 NUMERIC "1"
-- Retrieval info: PRIVATE: SCANOUTA NUMERIC "0"
-- Retrieval info: PRIVATE: SCANOUTB NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SHIFTOUTA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SHIFTOUTA_REG STRING "0"
-- Retrieval info: PRIVATE: SIGNA STRING "Signed"
-- Retrieval info: PRIVATE: SIGNA_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNA_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNA_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: SIGNA_REG STRING "0"
-- Retrieval info: PRIVATE: SIGNB STRING "Signed"
-- Retrieval info: PRIVATE: SIGNB_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_ACLR_SRC NUMERIC "3"
-- Retrieval info: PRIVATE: SIGNB_PIPE_CLK_SRC NUMERIC "0"
-- Retrieval info: PRIVATE: SIGNB_PIPE_REG STRING "0"
-- Retrieval info: PRIVATE: SIGNB_REG STRING "0"
-- Retrieval info: PRIVATE: SRCA0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SRCB0 STRING "Multiplier input"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: WIDTHA STRING "16"
-- Retrieval info: PRIVATE: WIDTHB STRING "16"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_PIPELINE_REGISTER1 STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: ADDNSUB_MULTIPLIER_REGISTER1 STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: DEDICATED_MULTIPLIER_CIRCUITRY STRING "AUTO"
-- Retrieval info: CONSTANT: INPUT_REGISTER_A0 STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: INPUT_REGISTER_B0 STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: INPUT_SOURCE_A0 STRING "DATAA"
-- Retrieval info: CONSTANT: INPUT_SOURCE_B0 STRING "DATAB"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altmult_add"
-- Retrieval info: CONSTANT: MULTIPLIER1_DIRECTION STRING "ADD"
-- Retrieval info: CONSTANT: MULTIPLIER_REGISTER0 STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: NUMBER_OF_MULTIPLIERS NUMERIC "1"
-- Retrieval info: CONSTANT: OUTPUT_REGISTER STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: PORT_ADDNSUB1 STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNA STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: PORT_SIGNB STRING "PORT_UNUSED"
-- Retrieval info: CONSTANT: REPRESENTATION_A STRING "SIGNED"
-- Retrieval info: CONSTANT: REPRESENTATION_B STRING "SIGNED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: SIGNED_PIPELINE_REGISTER_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: SIGNED_REGISTER_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: WIDTH_A NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_B NUMERIC "16"
-- Retrieval info: CONSTANT: WIDTH_RESULT NUMERIC "16"
-- Retrieval info: USED_PORT: dataa_0 0 0 16 0 INPUT GND "dataa_0[15..0]"
-- Retrieval info: USED_PORT: datab_0 0 0 16 0 INPUT GND "datab_0[15..0]"
-- Retrieval info: USED_PORT: result 0 0 16 0 OUTPUT GND "result[15..0]"
-- Retrieval info: CONNECT: result 0 0 16 0 @result 0 0 16 0
-- Retrieval info: CONNECT: @dataa 0 0 16 0 dataa_0 0 0 16 0
-- Retrieval info: CONNECT: @datab 0 0 16 0 datab_0 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL altmult_add0.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altmult_add0.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altmult_add0.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altmult_add0.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL altmult_add0_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
